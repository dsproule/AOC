module aoc4_tb;

endmodule