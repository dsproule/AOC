module aoc4_tb;

    logic clock, reset, write_en, read_en, ack, busy;
    logic [`BANK_ADDR_WIDTH-1:0] owner_row_addr;
    logic [`TX_DATA_WIDTH-1:0]   partial_vec_in, partial_vec_out;
    logic [`COL_ADDR_WIDTH-1:0]  col_addr;

    BankController dut (.*);

    initial forever #5 clock = ~clock;

    initial begin
        $dumpfile("aoc.vcd");
        $dumpvars(0, aoc4_tb);
    end

    task print_mem;
        for (int i = 0; i < `BANK_DEPTH; i++) begin
            $display("%0d: %1b", i, dut.bank.mem[i]);
        end
    endtask

    task write_mem(input logic [`TX_DATA_WIDTH-1:0]    partial_vec, 
                    input logic [`BANK_ADDR_WIDTH-1:0] row_i, 
                    input logic [`COL_ADDR_WIDTH-1:0]  col_i);
        @(negedge clock);
        write_en = 1'b1;
        partial_vec_in = partial_vec;
        owner_row_addr = row_i;
        col_addr = col_i;
        @(negedge clock);
        write_en = 1'b0;
        if (!ack) @(posedge ack);
        repeat (2) @(negedge clock);
    endtask

    int fd;
    int c;
    int done;

    int row_i, col_i;
    logic [`TX_DATA_WIDTH-1:0] partial_row_vec;

    initial begin
        fd = $fopen("input4.txt", "r");
        if (fd == 0) $fatal(1, "ERROR: Could not open input4.txt");

        clock    = 0;
        reset    = 1;
        read_en  = 0;
        write_en = 0;
        owner_row_addr = '0;
        partial_vec_in = '0;
        col_addr = 0;
        done     = 0;
        row_i    = 0;
        col_i    = 0;
        partial_row_vec = '0;

        repeat (3) @(negedge clock);
        reset = 0;

        // initialization of banks
        @(negedge clock);
        while (!done) begin
            c = $fgetc(fd);

            if (c == -1) begin
                done = 1;
            end else if (c == 10) begin
                write_mem(partial_row_vec, row_i, (`MAX_COLS / `TX_DATA_WIDTH) * `TX_DATA_WIDTH);
                col_i = 0;
                row_i++;
                
            end else begin
                if (col_i % `TX_DATA_WIDTH == 0 && col_i > 0) begin
                    write_mem(partial_row_vec, row_i, col_i - `TX_DATA_WIDTH);
                    partial_row_vec = '0;
                end
                partial_row_vec[col_i % `TX_DATA_WIDTH] = (c == "@");
                col_i++;
            end
        end

        print_mem;
        $finish;
    end

endmodule