`ifndef COMMON_SVH__
`define COMMON_SVH__

`define DATA_WIDTH 32

`endif